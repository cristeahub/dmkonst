library IEEE;
use IEEE.STD_LOGIC_1164.all;

package opcodes is

  constant FUNCTION_AND : std_logic_vector(3 downto 0) := "0000";

end opcodes;